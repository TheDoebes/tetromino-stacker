module tetrominos();
	// I/O
	
	// Internal Wiring
	reg tetromino[3:0][3:0][3:0];
	
	// Logic
	
	// Create Tetrominos
	assign tetromino[0][0] = {}
endmodule
		